library verilog;
use verilog.vl_types.all;
entity ram_test_vlg_vec_tst is
end ram_test_vlg_vec_tst;
